module nzp_module( input logic[15:0] data, input logic LD_CC, LD_BEN, input logic[2:0] currNZP,
						 output logic BEN );
endmodule
