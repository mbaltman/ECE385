module alu_module(input logic[15:0] A, B,input logic[1:0] s,  output logic[15:0] out);
endmodule
