module stateRegister(input logic [127:0] encoded_msg, mux_output, 
							input integer state_number, 
							input logic mux_enable);
							
endmodule 