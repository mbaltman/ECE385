/************************************************************************
Avalon-MM Interface for AES Decryption IP Core

Dong Kai Wang, Fall 2017

For use with ECE 385 Experiment 9
University of Illinois ECE Department

Register Map:

0-3 : 4x 32bit AES Key
4-7 : 4x 32bit AES Encrypted Message
8-11: 4x 32bit AES Decrypted Message
12: Not Used
13: Not Used
14: 32bit Start Register
15: 32bit Done Register

************************************************************************/

module avalon_aes_interface (
	// Avalon Clock Input
	input logic CLK,

	// Avalon Reset Input
	input logic RESET,

	// Avalon-MM Slave Signals
	input  logic AVL_READ,					// Avalon-MM Read
	input  logic AVL_WRITE,					// Avalon-MM Write
	input  logic AVL_CS,					// Avalon-MM Chip Select
	input  logic [3:0] AVL_BYTE_EN,			// Avalon-MM Byte Enable
	input  logic [3:0] AVL_ADDR,			// Avalon-MM Address
	input  logic [31:0] AVL_WRITEDATA,		// Avalon-MM Write Data
	output logic [31:0] AVL_READDATA,		// Avalon-MM Read Data

	// Exported Conduit
	output logic [31:0] EXPORT_DATA			// Exported Conduit Signal to LEDs
	);

	logic [31:0] registers [15:0];

	always_ff @ (posedge CLK) // write has 1 cycle of delay
	begin
		if (RESET)
		begin
			for (int i = 0; i < 16; i++)
			begin
				register_file[i] <= 32'b0; // clear everything to 0
			end
		end
		else if (AVL_WRITE && AVL_CS)
		begin
			register_file[AVL_ADDR][31:0] <= AVL_WRITEDATA[31:0]; // write data into corresponding address
		end
		else
		begin
			for (int i = 0; i < 16; i++)
			begin
				register_file[i] <= register_file[i]; // do nothing
			end
		end
	end

	always_comb // read has no delay
	begin
		if (AVL_READ && AVL_CS)
		begin
			AVL_READDATA[31:0] = register_file[AVL_ADDR][31:0]; // reading data out
		end
		else
		begin
			AVL_READDATA[31:0] = 32'b0; // not reading, high impedence
		end
	end

	assign EXPORT_DATA = {registers[0][31:16], registers[3][15:0]};

endmodule
